library verilog;
use verilog.vl_types.all;
entity seven_stage_monitor_vlg_vec_tst is
end seven_stage_monitor_vlg_vec_tst;
