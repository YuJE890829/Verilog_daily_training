library verilog;
use verilog.vl_types.all;
entity MUL4_vlg_vec_tst is
end MUL4_vlg_vec_tst;
