library verilog;
use verilog.vl_types.all;
entity D_flipflop_vlg_vec_tst is
end D_flipflop_vlg_vec_tst;
