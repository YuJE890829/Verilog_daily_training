library verilog;
use verilog.vl_types.all;
entity fourbits_CLGadder_vlg_vec_tst is
end fourbits_CLGadder_vlg_vec_tst;
