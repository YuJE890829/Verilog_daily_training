library verilog;
use verilog.vl_types.all;
entity ADDS4_vlg_vec_tst is
end ADDS4_vlg_vec_tst;
