library verilog;
use verilog.vl_types.all;
entity fourbits_adder_vlg_vec_tst is
end fourbits_adder_vlg_vec_tst;
