library verilog;
use verilog.vl_types.all;
entity priority_8bit_encoder_vlg_vec_tst is
end priority_8bit_encoder_vlg_vec_tst;
